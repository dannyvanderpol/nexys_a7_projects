----------------------------------------------------------------------------------------------------
-- Template
----------------------------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;

entity template is
    port(
        CLK_ : in std_logic
    );
end entity;


architecture behavior of template is
    

begin
    TEMPLATE : process (CLK_)
    begin
    
    end process;

end architecture;
